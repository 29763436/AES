library verilog;
use verilog.vl_types.all;
entity AESK_vlg_vec_tst is
end AESK_vlg_vec_tst;
